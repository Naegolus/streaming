-- megafunction wizard: %ALTREMOTE_UPDATE%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altremote_update 

-- ============================================================
-- File Name: altremote.vhd
-- Megafunction Name(s):
-- 			altremote_update
--
-- Simulation Library Files(s):
-- 			cycloneive;lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 10.1 Build 153 11/29/2010 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2010 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altremote_update CBX_AUTO_BLACKBOX="ALL" check_app_pof="false" DEVICE_FAMILY="Cyclone IV E" in_data_width=22 operation_mode="remote" out_data_width=29 busy clock data_in data_out param read_param read_source reconfig reset reset_timer write_param
--VERSION_BEGIN 10.1 cbx_altremote_update 2010:11:29:22:18:02:SJ cbx_cycloneii 2010:11:29:22:18:02:SJ cbx_lpm_add_sub 2010:11:29:22:18:02:SJ cbx_lpm_compare 2010:11:29:22:18:02:SJ cbx_lpm_counter 2010:11:29:22:18:02:SJ cbx_lpm_decode 2010:11:29:22:18:02:SJ cbx_lpm_shiftreg 2010:11:29:22:18:02:SJ cbx_mgl 2010:11:29:22:19:52:SJ cbx_stratix 2010:11:29:22:18:02:SJ cbx_stratixii 2010:11:29:22:18:02:SJ  VERSION_END

 LIBRARY cycloneive;
 USE cycloneive.all;

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = cycloneive_rublock 1 lpm_counter 2 reg 61 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  altremote_rmtupdt_51n IS 
	 PORT 
	 ( 
		 busy	:	OUT  STD_LOGIC;
		 clock	:	IN  STD_LOGIC;
		 data_in	:	IN  STD_LOGIC_VECTOR (21 DOWNTO 0) := (OTHERS => '0');
		 data_out	:	OUT  STD_LOGIC_VECTOR (28 DOWNTO 0);
		 param	:	IN  STD_LOGIC_VECTOR (2 DOWNTO 0) := (OTHERS => '0');
		 read_param	:	IN  STD_LOGIC := '0';
		 read_source	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0) := (OTHERS => '0');
		 reconfig	:	IN  STD_LOGIC := '0';
		 reset	:	IN  STD_LOGIC;
		 reset_timer	:	IN  STD_LOGIC := '0';
		 write_param	:	IN  STD_LOGIC := '0'
	 ); 
 END altremote_rmtupdt_51n;

 ARCHITECTURE RTL OF altremote_rmtupdt_51n IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "suppress_da_rule_internal=c104;suppress_da_rule_internal=C101;suppress_da_rule_internal=C103";

	 SIGNAL	 dffe10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe16	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe17	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe18	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe19	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe1a0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe1a1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_dffe1a_ena	:	STD_LOGIC_VECTOR(1 DOWNTO 0);
	 SIGNAL	 dffe20	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe22	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe23	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe24	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe25a	:	STD_LOGIC_VECTOR(6 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_dffe25a_ena	:	STD_LOGIC_VECTOR(6 DOWNTO 0);
	 SIGNAL	 dffe2a0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe2a1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe2a2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_dffe2a_ena	:	STD_LOGIC_VECTOR(2 DOWNTO 0);
	 SIGNAL	 dffe3a0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe3a1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe3a2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_dffe3a_ena	:	STD_LOGIC_VECTOR(2 DOWNTO 0);
	 SIGNAL	 dffe7a	:	STD_LOGIC_VECTOR(28 DOWNTO 0)
	 -- synopsys translate_off
	  := "00000000000000000000000000000"
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_dffe7a_clrn	:	STD_LOGIC_VECTOR(28 DOWNTO 0);
	 SIGNAL	 wire_dffe7a_ena	:	STD_LOGIC_VECTOR(28 DOWNTO 0);
	 SIGNAL	 dffe8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_cntr5_w_lg_w_q_range30w33w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cntr5_w_lg_w_q_range31w32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cntr5_q	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_cntr5_w_q_range30w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cntr5_w_q_range31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cntr6_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_sd4_regout	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w801w804w807w810w812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w801w804w840w841w842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w801w821w822w823w824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w815w816w817w818w819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w815w816w817w885w886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w815w816w844w845w846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w815w849w850w851w852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w815w849w907w908w909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w826w827w875w876w877w878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w826w827w828w829w830w831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w826w827w828w899w900w901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w826w888w889w890w891w892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w826w888w911w912w913w914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w868w869w870w871w873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w868w894w895w896w897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w834w880w881w882w883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w834w835w836w837w838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w834w835w903w904w905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w854w862w863w864w865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w854w855w856w857w858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w798w801w804w807w810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w798w801w804w840w841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w798w801w821w822w823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w798w815w816w817w818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w798w815w816w817w885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w798w815w816w844w845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w798w815w849w850w851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w798w815w849w907w908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w826w827w875w876w877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w826w827w828w829w830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w826w827w828w899w900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w826w888w889w890w891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w826w888w911w912w913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w868w869w870w871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w868w894w895w896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w834w880w881w882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w834w835w836w837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w834w835w903w904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w854w862w863w864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w854w855w856w857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w798w801w804w807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w798w801w804w840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w798w801w821w822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w798w815w816w817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w798w815w816w844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w798w815w849w850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w798w815w849w907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w826w827w875w876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w826w827w828w829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w826w827w828w899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w826w888w889w890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w826w888w911w912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w868w869w870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w868w894w895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w834w880w881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w834w835w836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w834w835w903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w854w862w863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w854w855w856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w798w801w804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w798w801w821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w798w815w816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w798w815w849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w826w827w875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w826w827w828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w826w888w889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w826w888w911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w868w869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w868w894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w834w880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w834w835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w854w862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w854w855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w798w801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w798w815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w826w827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w826w888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_idle949w950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_rsource_load5w6w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_rsource_load5w13w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_rsource_load5w17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_rsource_load5w23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_rsource_load5w27w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable93w96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable93w132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable93w136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable93w140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable93w144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable93w148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable93w152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable93w156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable93w160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable93w164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable93w168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable93w100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable93w172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable93w176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable93w180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable93w104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable93w108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable93w112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable93w116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable93w120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable93w124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable93w128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_source_update1007w1008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_data966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_init_counter962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_post972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_pre_data961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rsource_load7w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rsource_load14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rsource_load18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rsource_load24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rsource_load28w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rublock_regout_reg1013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_data984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_init_counter981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_post_data990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_pre_data980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range794w867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range794w833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_read_source_range1034w1035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_read_source_range1038w1039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_clear91w92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bit_counter_all_done983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bit_counter_param_start_match960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_data925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_init929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_init_counter927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_param948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_post924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_pre_data926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_source_update928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rsource_load5w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rsource_update_done957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_select_shift_nloop1012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_width_counter_all_done964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_width_counter_param_width_match965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_data919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_init923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_init_counter922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_load917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_param947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_post_data918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_pre_data920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_source_update921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_wait916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_wsource_update_done977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range794w795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range796w797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range799w800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range802w803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range805w806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range808w809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range811w872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_idle949w950w951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_read_source_range1034w1035w1036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_read_source_range1038w1039w1040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_source_update1007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rsource_load9w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rsource_load1w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_clear91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  bit_counter_all_done :	STD_LOGIC;
	 SIGNAL  bit_counter_clear :	STD_LOGIC;
	 SIGNAL  bit_counter_enable :	STD_LOGIC;
	 SIGNAL  bit_counter_param_start :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  bit_counter_param_start_match :	STD_LOGIC;
	 SIGNAL  combine_port :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  global_gnd :	STD_LOGIC;
	 SIGNAL  global_vcc :	STD_LOGIC;
	 SIGNAL  idle :	STD_LOGIC;
	 SIGNAL  param_decoder_param_latch :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  param_decoder_select :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  power_up :	STD_LOGIC;
	 SIGNAL  read_data :	STD_LOGIC;
	 SIGNAL  read_init :	STD_LOGIC;
	 SIGNAL  read_init_counter :	STD_LOGIC;
	 SIGNAL  read_post :	STD_LOGIC;
	 SIGNAL  read_pre_data :	STD_LOGIC;
	 SIGNAL  read_source_update :	STD_LOGIC;
	 SIGNAL  rsource_load :	STD_LOGIC;
	 SIGNAL  rsource_parallel_in :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  rsource_serial_out :	STD_LOGIC;
	 SIGNAL  rsource_shift_enable :	STD_LOGIC;
	 SIGNAL  rsource_state_par_ini :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rsource_update_done :	STD_LOGIC;
	 SIGNAL  rublock_captnupdt :	STD_LOGIC;
	 SIGNAL  rublock_clock :	STD_LOGIC;
	 SIGNAL  rublock_reconfig :	STD_LOGIC;
	 SIGNAL  rublock_reconfig_st :	STD_LOGIC;
	 SIGNAL  rublock_regin :	STD_LOGIC;
	 SIGNAL  rublock_regout :	STD_LOGIC;
	 SIGNAL  rublock_regout_reg :	STD_LOGIC;
	 SIGNAL  rublock_shiftnld :	STD_LOGIC;
	 SIGNAL  select_shift_nloop :	STD_LOGIC;
	 SIGNAL  shift_reg_clear :	STD_LOGIC;
	 SIGNAL  shift_reg_load_enable :	STD_LOGIC;
	 SIGNAL  shift_reg_serial_in :	STD_LOGIC;
	 SIGNAL  shift_reg_serial_out :	STD_LOGIC;
	 SIGNAL  shift_reg_shift_enable :	STD_LOGIC;
	 SIGNAL  start_bit_decoder_out :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  start_bit_decoder_param_select :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  w44w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  w74w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  width_counter_all_done :	STD_LOGIC;
	 SIGNAL  width_counter_clear :	STD_LOGIC;
	 SIGNAL  width_counter_enable :	STD_LOGIC;
	 SIGNAL  width_counter_param_width :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  width_counter_param_width_match :	STD_LOGIC;
	 SIGNAL  width_decoder_out :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  width_decoder_param_select :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  write_data :	STD_LOGIC;
	 SIGNAL  write_init :	STD_LOGIC;
	 SIGNAL  write_init_counter :	STD_LOGIC;
	 SIGNAL  write_load :	STD_LOGIC;
	 SIGNAL  write_post_data :	STD_LOGIC;
	 SIGNAL  write_pre_data :	STD_LOGIC;
	 SIGNAL  write_source_update :	STD_LOGIC;
	 SIGNAL  write_wait :	STD_LOGIC;
	 SIGNAL  wsource_state_par_ini :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wsource_update_done :	STD_LOGIC;
	 SIGNAL  wire_w_data_in_range95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_read_source_range1034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_read_source_range1038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rsource_parallel_in_range4w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rsource_state_par_ini_range12w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rsource_state_par_ini_range16w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_wsource_state_par_ini_range22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_wsource_state_par_ini_range26w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  cycloneive_rublock
	 PORT
	 ( 
		captnupdt	:	IN STD_LOGIC;
		clk	:	IN STD_LOGIC;
		rconfig	:	IN STD_LOGIC;
		regin	:	IN STD_LOGIC;
		regout	:	OUT STD_LOGIC;
		rsttimer	:	IN STD_LOGIC;
		shiftnld	:	IN STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w801w804w807w810w812w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w798w801w804w807w810w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w801w804w840w841w842w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w798w801w804w840w841w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w801w821w822w823w824w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w798w801w821w822w823w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w815w816w817w818w819w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w798w815w816w817w818w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w815w816w817w885w886w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w798w815w816w817w885w(0) AND wire_w_lg_w_param_decoder_param_latch_range811w872w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w815w816w844w845w846w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w798w815w816w844w845w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w815w849w850w851w852w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w798w815w849w850w851w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w815w849w907w908w909w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w798w815w849w907w908w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w826w827w875w876w877w878w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w826w827w875w876w877w(0) AND wire_w_lg_w_param_decoder_param_latch_range811w872w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w826w827w828w829w830w831w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w826w827w828w829w830w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w826w827w828w899w900w901w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w826w827w828w899w900w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w826w888w889w890w891w892w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w826w888w889w890w891w(0) AND wire_w_lg_w_param_decoder_param_latch_range811w872w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w826w888w911w912w913w914w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w826w888w911w912w913w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w868w869w870w871w873w(0) <= wire_w_lg_w_lg_w_lg_w868w869w870w871w(0) AND wire_w_lg_w_param_decoder_param_latch_range811w872w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w868w894w895w896w897w(0) <= wire_w_lg_w_lg_w_lg_w868w894w895w896w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w834w880w881w882w883w(0) <= wire_w_lg_w_lg_w_lg_w834w880w881w882w(0) AND wire_w_lg_w_param_decoder_param_latch_range811w872w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w834w835w836w837w838w(0) <= wire_w_lg_w_lg_w_lg_w834w835w836w837w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w834w835w903w904w905w(0) <= wire_w_lg_w_lg_w_lg_w834w835w903w904w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w854w862w863w864w865w(0) <= wire_w_lg_w_lg_w_lg_w854w862w863w864w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w854w855w856w857w858w(0) <= wire_w_lg_w_lg_w_lg_w854w855w856w857w(0) AND wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w798w801w804w807w810w(0) <= wire_w_lg_w_lg_w_lg_w798w801w804w807w(0) AND wire_w_lg_w_param_decoder_param_latch_range808w809w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w798w801w804w840w841w(0) <= wire_w_lg_w_lg_w_lg_w798w801w804w840w(0) AND wire_w_lg_w_param_decoder_param_latch_range808w809w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w798w801w821w822w823w(0) <= wire_w_lg_w_lg_w_lg_w798w801w821w822w(0) AND wire_w_lg_w_param_decoder_param_latch_range808w809w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w798w815w816w817w818w(0) <= wire_w_lg_w_lg_w_lg_w798w815w816w817w(0) AND wire_w_lg_w_param_decoder_param_latch_range808w809w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w798w815w816w817w885w(0) <= wire_w_lg_w_lg_w_lg_w798w815w816w817w(0) AND wire_w_param_decoder_param_latch_range808w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w798w815w816w844w845w(0) <= wire_w_lg_w_lg_w_lg_w798w815w816w844w(0) AND wire_w_lg_w_param_decoder_param_latch_range808w809w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w798w815w849w850w851w(0) <= wire_w_lg_w_lg_w_lg_w798w815w849w850w(0) AND wire_w_lg_w_param_decoder_param_latch_range808w809w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w798w815w849w907w908w(0) <= wire_w_lg_w_lg_w_lg_w798w815w849w907w(0) AND wire_w_lg_w_param_decoder_param_latch_range808w809w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w826w827w875w876w877w(0) <= wire_w_lg_w_lg_w_lg_w826w827w875w876w(0) AND wire_w_param_decoder_param_latch_range808w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w826w827w828w829w830w(0) <= wire_w_lg_w_lg_w_lg_w826w827w828w829w(0) AND wire_w_lg_w_param_decoder_param_latch_range808w809w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w826w827w828w899w900w(0) <= wire_w_lg_w_lg_w_lg_w826w827w828w899w(0) AND wire_w_lg_w_param_decoder_param_latch_range808w809w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w826w888w889w890w891w(0) <= wire_w_lg_w_lg_w_lg_w826w888w889w890w(0) AND wire_w_param_decoder_param_latch_range808w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w826w888w911w912w913w(0) <= wire_w_lg_w_lg_w_lg_w826w888w911w912w(0) AND wire_w_lg_w_param_decoder_param_latch_range808w809w(0);
	wire_w_lg_w_lg_w_lg_w868w869w870w871w(0) <= wire_w_lg_w_lg_w868w869w870w(0) AND wire_w_param_decoder_param_latch_range808w(0);
	wire_w_lg_w_lg_w_lg_w868w894w895w896w(0) <= wire_w_lg_w_lg_w868w894w895w(0) AND wire_w_lg_w_param_decoder_param_latch_range808w809w(0);
	wire_w_lg_w_lg_w_lg_w834w880w881w882w(0) <= wire_w_lg_w_lg_w834w880w881w(0) AND wire_w_param_decoder_param_latch_range808w(0);
	wire_w_lg_w_lg_w_lg_w834w835w836w837w(0) <= wire_w_lg_w_lg_w834w835w836w(0) AND wire_w_lg_w_param_decoder_param_latch_range808w809w(0);
	wire_w_lg_w_lg_w_lg_w834w835w903w904w(0) <= wire_w_lg_w_lg_w834w835w903w(0) AND wire_w_lg_w_param_decoder_param_latch_range808w809w(0);
	wire_w_lg_w_lg_w_lg_w854w862w863w864w(0) <= wire_w_lg_w_lg_w854w862w863w(0) AND wire_w_lg_w_param_decoder_param_latch_range808w809w(0);
	wire_w_lg_w_lg_w_lg_w854w855w856w857w(0) <= wire_w_lg_w_lg_w854w855w856w(0) AND wire_w_lg_w_param_decoder_param_latch_range808w809w(0);
	wire_w_lg_w_lg_w_lg_w798w801w804w807w(0) <= wire_w_lg_w_lg_w798w801w804w(0) AND wire_w_lg_w_param_decoder_param_latch_range805w806w(0);
	wire_w_lg_w_lg_w_lg_w798w801w804w840w(0) <= wire_w_lg_w_lg_w798w801w804w(0) AND wire_w_param_decoder_param_latch_range805w(0);
	wire_w_lg_w_lg_w_lg_w798w801w821w822w(0) <= wire_w_lg_w_lg_w798w801w821w(0) AND wire_w_lg_w_param_decoder_param_latch_range805w806w(0);
	wire_w_lg_w_lg_w_lg_w798w815w816w817w(0) <= wire_w_lg_w_lg_w798w815w816w(0) AND wire_w_lg_w_param_decoder_param_latch_range805w806w(0);
	wire_w_lg_w_lg_w_lg_w798w815w816w844w(0) <= wire_w_lg_w_lg_w798w815w816w(0) AND wire_w_param_decoder_param_latch_range805w(0);
	wire_w_lg_w_lg_w_lg_w798w815w849w850w(0) <= wire_w_lg_w_lg_w798w815w849w(0) AND wire_w_lg_w_param_decoder_param_latch_range805w806w(0);
	wire_w_lg_w_lg_w_lg_w798w815w849w907w(0) <= wire_w_lg_w_lg_w798w815w849w(0) AND wire_w_param_decoder_param_latch_range805w(0);
	wire_w_lg_w_lg_w_lg_w826w827w875w876w(0) <= wire_w_lg_w_lg_w826w827w875w(0) AND wire_w_lg_w_param_decoder_param_latch_range805w806w(0);
	wire_w_lg_w_lg_w_lg_w826w827w828w829w(0) <= wire_w_lg_w_lg_w826w827w828w(0) AND wire_w_lg_w_param_decoder_param_latch_range805w806w(0);
	wire_w_lg_w_lg_w_lg_w826w827w828w899w(0) <= wire_w_lg_w_lg_w826w827w828w(0) AND wire_w_param_decoder_param_latch_range805w(0);
	wire_w_lg_w_lg_w_lg_w826w888w889w890w(0) <= wire_w_lg_w_lg_w826w888w889w(0) AND wire_w_lg_w_param_decoder_param_latch_range805w806w(0);
	wire_w_lg_w_lg_w_lg_w826w888w911w912w(0) <= wire_w_lg_w_lg_w826w888w911w(0) AND wire_w_param_decoder_param_latch_range805w(0);
	wire_w_lg_w_lg_w868w869w870w(0) <= wire_w_lg_w868w869w(0) AND wire_w_lg_w_param_decoder_param_latch_range805w806w(0);
	wire_w_lg_w_lg_w868w894w895w(0) <= wire_w_lg_w868w894w(0) AND wire_w_param_decoder_param_latch_range805w(0);
	wire_w_lg_w_lg_w834w880w881w(0) <= wire_w_lg_w834w880w(0) AND wire_w_lg_w_param_decoder_param_latch_range805w806w(0);
	wire_w_lg_w_lg_w834w835w836w(0) <= wire_w_lg_w834w835w(0) AND wire_w_lg_w_param_decoder_param_latch_range805w806w(0);
	wire_w_lg_w_lg_w834w835w903w(0) <= wire_w_lg_w834w835w(0) AND wire_w_param_decoder_param_latch_range805w(0);
	wire_w_lg_w_lg_w854w862w863w(0) <= wire_w_lg_w854w862w(0) AND wire_w_param_decoder_param_latch_range805w(0);
	wire_w_lg_w_lg_w854w855w856w(0) <= wire_w_lg_w854w855w(0) AND wire_w_lg_w_param_decoder_param_latch_range805w806w(0);
	wire_w_lg_w_lg_w798w801w804w(0) <= wire_w_lg_w798w801w(0) AND wire_w_lg_w_param_decoder_param_latch_range802w803w(0);
	wire_w_lg_w_lg_w798w801w821w(0) <= wire_w_lg_w798w801w(0) AND wire_w_param_decoder_param_latch_range802w(0);
	wire_w_lg_w_lg_w798w815w816w(0) <= wire_w_lg_w798w815w(0) AND wire_w_lg_w_param_decoder_param_latch_range802w803w(0);
	wire_w_lg_w_lg_w798w815w849w(0) <= wire_w_lg_w798w815w(0) AND wire_w_param_decoder_param_latch_range802w(0);
	wire_w_lg_w_lg_w826w827w875w(0) <= wire_w_lg_w826w827w(0) AND wire_w_lg_w_param_decoder_param_latch_range802w803w(0);
	wire_w_lg_w_lg_w826w827w828w(0) <= wire_w_lg_w826w827w(0) AND wire_w_param_decoder_param_latch_range802w(0);
	wire_w_lg_w_lg_w826w888w889w(0) <= wire_w_lg_w826w888w(0) AND wire_w_lg_w_param_decoder_param_latch_range802w803w(0);
	wire_w_lg_w_lg_w826w888w911w(0) <= wire_w_lg_w826w888w(0) AND wire_w_param_decoder_param_latch_range802w(0);
	wire_w_lg_w868w869w(0) <= wire_w868w(0) AND wire_w_lg_w_param_decoder_param_latch_range802w803w(0);
	wire_w_lg_w868w894w(0) <= wire_w868w(0) AND wire_w_param_decoder_param_latch_range802w(0);
	wire_w_lg_w834w880w(0) <= wire_w834w(0) AND wire_w_lg_w_param_decoder_param_latch_range802w803w(0);
	wire_w_lg_w834w835w(0) <= wire_w834w(0) AND wire_w_param_decoder_param_latch_range802w(0);
	wire_w_lg_w854w862w(0) <= wire_w854w(0) AND wire_w_lg_w_param_decoder_param_latch_range802w803w(0);
	wire_w_lg_w854w855w(0) <= wire_w854w(0) AND wire_w_param_decoder_param_latch_range802w(0);
	wire_w_lg_w798w801w(0) <= wire_w798w(0) AND wire_w_lg_w_param_decoder_param_latch_range799w800w(0);
	wire_w_lg_w798w815w(0) <= wire_w798w(0) AND wire_w_param_decoder_param_latch_range799w(0);
	wire_w_lg_w826w827w(0) <= wire_w826w(0) AND wire_w_lg_w_param_decoder_param_latch_range799w800w(0);
	wire_w_lg_w826w888w(0) <= wire_w826w(0) AND wire_w_param_decoder_param_latch_range799w(0);
	wire_w_lg_w_lg_idle949w950w(0) <= wire_w_lg_idle949w(0) AND wire_w_lg_write_param947w(0);
	wire_w868w(0) <= wire_w_lg_w_param_decoder_param_latch_range794w867w(0) AND wire_w_lg_w_param_decoder_param_latch_range799w800w(0);
	wire_w834w(0) <= wire_w_lg_w_param_decoder_param_latch_range794w833w(0) AND wire_w_lg_w_param_decoder_param_latch_range799w800w(0);
	wire_w854w(0) <= wire_w_lg_w_param_decoder_param_latch_range794w833w(0) AND wire_w_param_decoder_param_latch_range799w(0);
	wire_w_lg_w_lg_rsource_load5w6w(0) <= wire_w_lg_rsource_load5w(0) AND dffe1a1;
	wire_w_lg_w_lg_rsource_load5w13w(0) <= wire_w_lg_rsource_load5w(0) AND dffe2a1;
	wire_w_lg_w_lg_rsource_load5w17w(0) <= wire_w_lg_rsource_load5w(0) AND dffe2a2;
	wire_w_lg_w_lg_rsource_load5w23w(0) <= wire_w_lg_rsource_load5w(0) AND dffe3a1;
	wire_w_lg_w_lg_rsource_load5w27w(0) <= wire_w_lg_rsource_load5w(0) AND dffe3a2;
	wire_w_lg_w_lg_shift_reg_load_enable93w96w(0) <= wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(1);
	wire_w_lg_w_lg_shift_reg_load_enable93w132w(0) <= wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(10);
	wire_w_lg_w_lg_shift_reg_load_enable93w136w(0) <= wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(11);
	wire_w_lg_w_lg_shift_reg_load_enable93w140w(0) <= wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(12);
	wire_w_lg_w_lg_shift_reg_load_enable93w144w(0) <= wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(13);
	wire_w_lg_w_lg_shift_reg_load_enable93w148w(0) <= wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(14);
	wire_w_lg_w_lg_shift_reg_load_enable93w152w(0) <= wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(15);
	wire_w_lg_w_lg_shift_reg_load_enable93w156w(0) <= wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(16);
	wire_w_lg_w_lg_shift_reg_load_enable93w160w(0) <= wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(17);
	wire_w_lg_w_lg_shift_reg_load_enable93w164w(0) <= wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(18);
	wire_w_lg_w_lg_shift_reg_load_enable93w168w(0) <= wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(19);
	wire_w_lg_w_lg_shift_reg_load_enable93w100w(0) <= wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(2);
	wire_w_lg_w_lg_shift_reg_load_enable93w172w(0) <= wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(20);
	wire_w_lg_w_lg_shift_reg_load_enable93w176w(0) <= wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(21);
	wire_w_lg_w_lg_shift_reg_load_enable93w180w(0) <= wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(22);
	wire_w_lg_w_lg_shift_reg_load_enable93w104w(0) <= wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(3);
	wire_w_lg_w_lg_shift_reg_load_enable93w108w(0) <= wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(4);
	wire_w_lg_w_lg_shift_reg_load_enable93w112w(0) <= wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(5);
	wire_w_lg_w_lg_shift_reg_load_enable93w116w(0) <= wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(6);
	wire_w_lg_w_lg_shift_reg_load_enable93w120w(0) <= wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(7);
	wire_w_lg_w_lg_shift_reg_load_enable93w124w(0) <= wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(8);
	wire_w_lg_w_lg_shift_reg_load_enable93w128w(0) <= wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(9);
	wire_w798w(0) <= wire_w_lg_w_param_decoder_param_latch_range794w795w(0) AND wire_w_lg_w_param_decoder_param_latch_range796w797w(0);
	wire_w826w(0) <= wire_w_lg_w_param_decoder_param_latch_range794w795w(0) AND wire_w_param_decoder_param_latch_range796w(0);
	wire_w_lg_w_lg_read_source_update1007w1008w(0) <= wire_w_lg_read_source_update1007w(0) AND rsource_serial_out;
	wire_w_lg_idle949w(0) <= idle AND wire_w_lg_read_param948w(0);
	wire_w_lg_read_data966w(0) <= read_data AND wire_w_lg_width_counter_param_width_match965w(0);
	wire_w_lg_read_init_counter962w(0) <= read_init_counter AND wire_w_lg_bit_counter_param_start_match960w(0);
	wire_w_lg_read_post972w(0) <= read_post AND wire_w_lg_width_counter_all_done964w(0);
	wire_w_lg_read_pre_data961w(0) <= read_pre_data AND wire_w_lg_bit_counter_param_start_match960w(0);
	wire_w_lg_rsource_load7w(0) <= rsource_load AND wire_w_rsource_parallel_in_range4w(0);
	wire_w_lg_rsource_load14w(0) <= rsource_load AND wire_w_rsource_state_par_ini_range12w(0);
	wire_w_lg_rsource_load18w(0) <= rsource_load AND wire_w_rsource_state_par_ini_range16w(0);
	wire_w_lg_rsource_load24w(0) <= rsource_load AND wire_w_wsource_state_par_ini_range22w(0);
	wire_w_lg_rsource_load28w(0) <= rsource_load AND wire_w_wsource_state_par_ini_range26w(0);
	wire_w_lg_rublock_regout_reg1013w(0) <= rublock_regout_reg AND wire_w_lg_select_shift_nloop1012w(0);
	wire_w_lg_shift_reg_load_enable97w(0) <= shift_reg_load_enable AND wire_w_data_in_range95w(0);
	wire_w_lg_shift_reg_load_enable137w(0) <= shift_reg_load_enable AND wire_w_data_in_range135w(0);
	wire_w_lg_shift_reg_load_enable141w(0) <= shift_reg_load_enable AND wire_w_data_in_range139w(0);
	wire_w_lg_shift_reg_load_enable145w(0) <= shift_reg_load_enable AND wire_w_data_in_range143w(0);
	wire_w_lg_shift_reg_load_enable149w(0) <= shift_reg_load_enable AND wire_w_data_in_range147w(0);
	wire_w_lg_shift_reg_load_enable153w(0) <= shift_reg_load_enable AND wire_w_data_in_range151w(0);
	wire_w_lg_shift_reg_load_enable157w(0) <= shift_reg_load_enable AND wire_w_data_in_range155w(0);
	wire_w_lg_shift_reg_load_enable161w(0) <= shift_reg_load_enable AND wire_w_data_in_range159w(0);
	wire_w_lg_shift_reg_load_enable165w(0) <= shift_reg_load_enable AND wire_w_data_in_range163w(0);
	wire_w_lg_shift_reg_load_enable169w(0) <= shift_reg_load_enable AND wire_w_data_in_range167w(0);
	wire_w_lg_shift_reg_load_enable173w(0) <= shift_reg_load_enable AND wire_w_data_in_range171w(0);
	wire_w_lg_shift_reg_load_enable101w(0) <= shift_reg_load_enable AND wire_w_data_in_range99w(0);
	wire_w_lg_shift_reg_load_enable177w(0) <= shift_reg_load_enable AND wire_w_data_in_range175w(0);
	wire_w_lg_shift_reg_load_enable181w(0) <= shift_reg_load_enable AND wire_w_data_in_range179w(0);
	wire_w_lg_shift_reg_load_enable105w(0) <= shift_reg_load_enable AND wire_w_data_in_range103w(0);
	wire_w_lg_shift_reg_load_enable109w(0) <= shift_reg_load_enable AND wire_w_data_in_range107w(0);
	wire_w_lg_shift_reg_load_enable113w(0) <= shift_reg_load_enable AND wire_w_data_in_range111w(0);
	wire_w_lg_shift_reg_load_enable117w(0) <= shift_reg_load_enable AND wire_w_data_in_range115w(0);
	wire_w_lg_shift_reg_load_enable121w(0) <= shift_reg_load_enable AND wire_w_data_in_range119w(0);
	wire_w_lg_shift_reg_load_enable125w(0) <= shift_reg_load_enable AND wire_w_data_in_range123w(0);
	wire_w_lg_shift_reg_load_enable129w(0) <= shift_reg_load_enable AND wire_w_data_in_range127w(0);
	wire_w_lg_shift_reg_load_enable133w(0) <= shift_reg_load_enable AND wire_w_data_in_range131w(0);
	wire_w_lg_write_data984w(0) <= write_data AND wire_w_lg_width_counter_param_width_match965w(0);
	wire_w_lg_write_init_counter981w(0) <= write_init_counter AND wire_w_lg_bit_counter_param_start_match960w(0);
	wire_w_lg_write_post_data990w(0) <= write_post_data AND wire_w_lg_bit_counter_all_done983w(0);
	wire_w_lg_write_pre_data980w(0) <= write_pre_data AND wire_w_lg_bit_counter_param_start_match960w(0);
	wire_w_lg_w_param_decoder_param_latch_range794w867w(0) <= wire_w_param_decoder_param_latch_range794w(0) AND wire_w_lg_w_param_decoder_param_latch_range796w797w(0);
	wire_w_lg_w_param_decoder_param_latch_range794w833w(0) <= wire_w_param_decoder_param_latch_range794w(0) AND wire_w_param_decoder_param_latch_range796w(0);
	wire_w_lg_w_read_source_range1034w1035w(0) <= wire_w_read_source_range1034w(0) AND read_param;
	wire_w_lg_w_read_source_range1038w1039w(0) <= wire_w_read_source_range1038w(0) AND read_param;
	wire_w_lg_w_lg_shift_reg_clear91w92w(0) <= NOT wire_w_lg_shift_reg_clear91w(0);
	wire_w_lg_bit_counter_all_done983w(0) <= NOT bit_counter_all_done;
	wire_w_lg_bit_counter_param_start_match960w(0) <= NOT bit_counter_param_start_match;
	wire_w_lg_idle930w(0) <= NOT idle;
	wire_w_lg_read_data925w(0) <= NOT read_data;
	wire_w_lg_read_init929w(0) <= NOT read_init;
	wire_w_lg_read_init_counter927w(0) <= NOT read_init_counter;
	wire_w_lg_read_param948w(0) <= NOT read_param;
	wire_w_lg_read_post924w(0) <= NOT read_post;
	wire_w_lg_read_pre_data926w(0) <= NOT read_pre_data;
	wire_w_lg_read_source_update928w(0) <= NOT read_source_update;
	wire_w_lg_rsource_load5w(0) <= NOT rsource_load;
	wire_w_lg_rsource_update_done957w(0) <= NOT rsource_update_done;
	wire_w_lg_select_shift_nloop1012w(0) <= NOT select_shift_nloop;
	wire_w_lg_shift_reg_load_enable93w(0) <= NOT shift_reg_load_enable;
	wire_w_lg_width_counter_all_done964w(0) <= NOT width_counter_all_done;
	wire_w_lg_width_counter_param_width_match965w(0) <= NOT width_counter_param_width_match;
	wire_w_lg_write_data919w(0) <= NOT write_data;
	wire_w_lg_write_init923w(0) <= NOT write_init;
	wire_w_lg_write_init_counter922w(0) <= NOT write_init_counter;
	wire_w_lg_write_load917w(0) <= NOT write_load;
	wire_w_lg_write_param947w(0) <= NOT write_param;
	wire_w_lg_write_post_data918w(0) <= NOT write_post_data;
	wire_w_lg_write_pre_data920w(0) <= NOT write_pre_data;
	wire_w_lg_write_source_update921w(0) <= NOT write_source_update;
	wire_w_lg_write_wait916w(0) <= NOT write_wait;
	wire_w_lg_wsource_update_done977w(0) <= NOT wsource_update_done;
	wire_w_lg_w_param_decoder_param_latch_range794w795w(0) <= NOT wire_w_param_decoder_param_latch_range794w(0);
	wire_w_lg_w_param_decoder_param_latch_range796w797w(0) <= NOT wire_w_param_decoder_param_latch_range796w(0);
	wire_w_lg_w_param_decoder_param_latch_range799w800w(0) <= NOT wire_w_param_decoder_param_latch_range799w(0);
	wire_w_lg_w_param_decoder_param_latch_range802w803w(0) <= NOT wire_w_param_decoder_param_latch_range802w(0);
	wire_w_lg_w_param_decoder_param_latch_range805w806w(0) <= NOT wire_w_param_decoder_param_latch_range805w(0);
	wire_w_lg_w_param_decoder_param_latch_range808w809w(0) <= NOT wire_w_param_decoder_param_latch_range808w(0);
	wire_w_lg_w_param_decoder_param_latch_range811w872w(0) <= NOT wire_w_param_decoder_param_latch_range811w(0);
	wire_w_lg_w_lg_w_lg_idle949w950w951w(0) <= wire_w_lg_w_lg_idle949w950w(0) OR write_wait;
	wire_w_lg_w_lg_w_read_source_range1034w1035w1036w(0) <= wire_w_lg_w_read_source_range1034w1035w(0) OR write_param;
	wire_w_lg_w_lg_w_read_source_range1038w1039w1040w(0) <= wire_w_lg_w_read_source_range1038w1039w(0) OR write_param;
	wire_w_lg_read_source_update1007w(0) <= read_source_update OR write_source_update;
	wire_w_lg_rsource_load9w(0) <= rsource_load OR global_vcc;
	wire_w_lg_rsource_load1w(0) <= rsource_load OR rsource_shift_enable;
	wire_w_lg_shift_reg_clear91w(0) <= shift_reg_clear OR reset;
	wire_w_lg_shift_reg_load_enable90w(0) <= shift_reg_load_enable OR shift_reg_shift_enable;
	bit_counter_all_done <= ((((wire_cntr5_w_lg_w_q_range30w33w(0) AND (NOT wire_cntr5_q(2))) AND wire_cntr5_q(3)) AND (NOT wire_cntr5_q(4))) AND wire_cntr5_q(5));
	bit_counter_clear <= (rsource_update_done OR wsource_update_done);
	bit_counter_enable <= (((((((((rsource_update_done OR wsource_update_done) OR read_init_counter) OR write_init_counter) OR read_pre_data) OR write_pre_data) OR read_data) OR write_data) OR read_post) OR write_post_data);
	bit_counter_param_start <= start_bit_decoder_out;
	bit_counter_param_start_match <= ((((((NOT w44w(0)) AND (NOT w44w(1))) AND (NOT w44w(2))) AND (NOT w44w(3))) AND (NOT w44w(4))) AND (NOT w44w(5)));
	busy <= wire_w_lg_idle930w(0);
	combine_port <= ( read_param & write_param & read_source & param);
	data_out <= dffe7a;
	global_gnd <= '0';
	global_vcc <= '1';
	idle <= dffe8;
	param_decoder_param_latch <= dffe25a;
	param_decoder_select <= ( wire_w_lg_w_lg_w_lg_w_lg_w_lg_w826w888w911w912w913w914w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w815w849w907w908w909w & wire_w_lg_w_lg_w_lg_w_lg_w834w835w903w904w905w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w826w827w828w899w900w901w & wire_w_lg_w_lg_w_lg_w_lg_w868w894w895w896w897w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w826w888w889w890w891w892w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w815w816w817w885w886w & wire_w_lg_w_lg_w_lg_w_lg_w834w880w881w882w883w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w826w827w875w876w877w878w & wire_w_lg_w_lg_w_lg_w_lg_w868w869w870w871w873w & wire_w_lg_w_lg_w_lg_w_lg_w854w862w863w864w865w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w815w816w844w845w846w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w801w804w840w841w842w & wire_w_lg_w_lg_w_lg_w_lg_w854w855w856w857w858w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w815w849w850w851w852w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w801w821w822w823w824w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w815w816w844w845w846w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w801w804w840w841w842w & wire_w_lg_w_lg_w_lg_w_lg_w834w835w836w837w838w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w826w827w828w829w830w831w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w801w821w822w823w824w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w815w816w817w818w819w & wire_w_lg_w_lg_w_lg_w_lg_w_lg_w798w801w804w807w810w812w);
	power_up <= ((((((((((((((wire_w_lg_idle930w(0) AND wire_w_lg_read_init929w(0)) AND wire_w_lg_read_source_update928w(0)) AND wire_w_lg_read_init_counter927w(0)) AND wire_w_lg_read_pre_data926w(0)) AND wire_w_lg_read_data925w(0)) AND wire_w_lg_read_post924w(0)) AND wire_w_lg_write_init923w(0)) AND wire_w_lg_write_init_counter922w(0)) AND wire_w_lg_write_source_update921w(0)) AND wire_w_lg_write_pre_data920w(0)) AND wire_w_lg_write_data919w(0)) AND wire_w_lg_write_post_data918w(0)) AND wire_w_lg_write_load917w(0)) AND wire_w_lg_write_wait916w(0));
	read_data <= dffe14;
	read_init <= dffe10;
	read_init_counter <= dffe12;
	read_post <= dffe15;
	read_pre_data <= dffe13;
	read_source_update <= dffe11;
	rsource_load <= (idle AND (write_param OR read_param));
	rsource_parallel_in <= ( wire_w_lg_w_lg_w_read_source_range1038w1039w1040w & wire_w_lg_w_lg_w_read_source_range1034w1035w1036w);
	rsource_serial_out <= dffe1a0;
	rsource_shift_enable <= wire_w_lg_read_source_update1007w(0);
	rsource_state_par_ini <= ( read_param & global_gnd & global_gnd);
	rsource_update_done <= dffe2a0;
	rublock_captnupdt <= wire_w_lg_write_load917w(0);
	rublock_clock <= (NOT (clock OR dffe9));
	rublock_reconfig <= rublock_reconfig_st;
	rublock_reconfig_st <= (idle AND reconfig);
	rublock_regin <= ((((wire_w_lg_rublock_regout_reg1013w(0) AND wire_w_lg_read_source_update928w(0)) AND wire_w_lg_write_source_update921w(0)) OR (((shift_reg_serial_out AND select_shift_nloop) AND wire_w_lg_read_source_update928w(0)) AND wire_w_lg_write_source_update921w(0))) OR wire_w_lg_w_lg_read_source_update1007w1008w(0));
	rublock_regout <= wire_sd4_regout;
	rublock_regout_reg <= dffe24;
	rublock_shiftnld <= (((((((read_pre_data OR write_pre_data) OR read_data) OR write_data) OR read_post) OR write_post_data) OR read_source_update) OR write_source_update);
	select_shift_nloop <= (wire_w_lg_read_data966w(0) OR wire_w_lg_write_data984w(0));
	shift_reg_clear <= read_init;
	shift_reg_load_enable <= (idle AND write_param);
	shift_reg_serial_in <= (rublock_regout_reg AND select_shift_nloop);
	shift_reg_serial_out <= dffe7a(0);
	shift_reg_shift_enable <= (((read_data OR write_data) OR read_post) OR write_post_data);
	start_bit_decoder_out <= ((((((((((((((((((((((( "0" & start_bit_decoder_param_select(0) & start_bit_decoder_param_select(0) & start_bit_decoder_param_select(0) & start_bit_decoder_param_select(0) & "0") OR ( "0" & "0" & "0" & "0" & "0" & "0")) OR ( "0" & start_bit_decoder_param_select(2) & start_bit_decoder_param_select(2) & start_bit_decoder_param_select(2) & start_bit_decoder_param_select(2) & "0")) OR ( "0" & "0" & "0" & "0" & "0" & "0")) OR ( "0" & start_bit_decoder_param_select(4) & start_bit_decoder_param_select(4) & start_bit_decoder_param_select(4) & "0" & start_bit_decoder_param_select(4))) OR ( "0" & start_bit_decoder_param_select(5) & start_bit_decoder_param_select(5) & start_bit_decoder_param_select(5) & start_bit_decoder_param_select(5) & "0")) OR ( "0" & "0" & "0" & "0" & "0" & "0")) OR ( "0" & start_bit_decoder_param_select(7) & start_bit_decoder_param_select(7) & "0" & "0" & "0")) OR ( "0" & "0" & "0" & "0" & "0" & "0")) OR ( "0" & start_bit_decoder_param_select(9) & start_bit_decoder_param_select(9) & "0" & start_bit_decoder_param_select(9) & "0")) OR ( "0" & start_bit_decoder_param_select(10) & start_bit_decoder_param_select(10) & "0" & "0" & "0")) OR ( "0" & "0" & "0" & "0" & "0" & "0")) OR ( "0" & start_bit_decoder_param_select(12) & start_bit_decoder_param_select(12) & "0" & start_bit_decoder_param_select(12) & "0")) OR ( start_bit_decoder_param_select(13) & "0" & "0" & start_bit_decoder_param_select(13) & "0" & start_bit_decoder_param_select(13))) OR ( "0" & "0" & "0" & "0" & "0" & "0")) OR ( start_bit_decoder_param_select(15) & "0" & "0" & "0" & start_bit_decoder_param_select(15) & start_bit_decoder_param_select(15))) OR ( "0" & "0" & start_bit_decoder_param_select(16) & start_bit_decoder_param_select(16) & "0" & "0")) OR ( start_bit_decoder_param_select(17) & "0" & "0" & start_bit_decoder_param_select(17) & "0" & "0")) OR ( start_bit_decoder_param_select(18) & "0" & "0" & start_bit_decoder_param_select(18) & "0" & start_bit_decoder_param_select(18))) OR ( "0" & "0" & "0" & "0" & "0" & "0"
)) OR ( start_bit_decoder_param_select(20) & "0" & "0" & "0" & start_bit_decoder_param_select(20) & start_bit_decoder_param_select(20))) OR ( "0" & "0" & start_bit_decoder_param_select(21) & start_bit_decoder_param_select(21) & "0" & "0")) OR ( start_bit_decoder_param_select(22) & "0" & "0" & start_bit_decoder_param_select(22) & "0" & "0"));
	start_bit_decoder_param_select <= param_decoder_select;
	w44w <= (wire_cntr5_q XOR bit_counter_param_start);
	w74w <= (wire_cntr6_q XOR width_counter_param_width);
	width_counter_all_done <= (((((NOT wire_cntr6_q(0)) AND (NOT wire_cntr6_q(1))) AND wire_cntr6_q(2)) AND wire_cntr6_q(3)) AND wire_cntr6_q(4));
	width_counter_clear <= (rsource_update_done OR wsource_update_done);
	width_counter_enable <= ((read_data OR write_data) OR read_post);
	width_counter_param_width <= width_decoder_out;
	width_counter_param_width_match <= (((((NOT w74w(0)) AND (NOT w74w(1))) AND (NOT w74w(2))) AND (NOT w74w(3))) AND (NOT w74w(4)));
	width_decoder_out <= ((((((((((((((((((((((( "0" & "0" & "0" & width_decoder_param_select(0) & "0") OR ( width_decoder_param_select(1) & width_decoder_param_select(1) & "0" & "0" & "0")) OR ( "0" & "0" & "0" & width_decoder_param_select(2) & "0")) OR ( width_decoder_param_select(3) & width_decoder_param_select(3) & width_decoder_param_select(3) & "0" & width_decoder_param_select(3))) OR ( "0" & "0" & "0" & "0" & width_decoder_param_select(4))) OR ( "0" & "0" & "0" & width_decoder_param_select(5) & "0")) OR ( width_decoder_param_select(6) & width_decoder_param_select(6) & "0" & "0" & "0")) OR ( "0" & "0" & "0" & width_decoder_param_select(7) & "0")) OR ( width_decoder_param_select(8) & width_decoder_param_select(8) & "0" & "0" & "0")) OR ( "0" & "0" & width_decoder_param_select(9) & "0" & width_decoder_param_select(9))) OR ( "0" & "0" & "0" & width_decoder_param_select(10) & "0")) OR ( width_decoder_param_select(11) & width_decoder_param_select(11) & "0" & "0" & "0")) OR ( "0" & "0" & width_decoder_param_select(12) & "0" & width_decoder_param_select(12))) OR ( "0" & "0" & "0" & "0" & width_decoder_param_select(13))) OR ( "0" & width_decoder_param_select(14) & width_decoder_param_select(14) & "0" & "0")) OR ( "0" & "0" & "0" & "0" & width_decoder_param_select(15))) OR ( width_decoder_param_select(16) & "0" & width_decoder_param_select(16) & width_decoder_param_select(16) & "0")) OR ( "0" & "0" & "0" & "0" & width_decoder_param_select(17))) OR ( "0" & "0" & "0" & "0" & width_decoder_param_select(18))) OR ( "0" & width_decoder_param_select(19) & width_decoder_param_select(19) & "0" & "0")) OR ( "0" & "0" & "0" & "0" & width_decoder_param_select(20))) OR ( width_decoder_param_select(21) & "0" & width_decoder_param_select(21) & width_decoder_param_select(21) & "0")) OR ( "0" & "0" & "0" & "0" & width_decoder_param_select(22)));
	width_decoder_param_select <= param_decoder_select;
	write_data <= dffe20;
	write_init <= dffe16;
	write_init_counter <= dffe18;
	write_load <= dffe22;
	write_post_data <= dffe21;
	write_pre_data <= dffe19;
	write_source_update <= dffe17;
	write_wait <= dffe23;
	wsource_state_par_ini <= ( write_param & global_gnd & global_gnd);
	wsource_update_done <= dffe3a0;
	wire_w_data_in_range95w(0) <= data_in(0);
	wire_w_data_in_range135w(0) <= data_in(10);
	wire_w_data_in_range139w(0) <= data_in(11);
	wire_w_data_in_range143w(0) <= data_in(12);
	wire_w_data_in_range147w(0) <= data_in(13);
	wire_w_data_in_range151w(0) <= data_in(14);
	wire_w_data_in_range155w(0) <= data_in(15);
	wire_w_data_in_range159w(0) <= data_in(16);
	wire_w_data_in_range163w(0) <= data_in(17);
	wire_w_data_in_range167w(0) <= data_in(18);
	wire_w_data_in_range171w(0) <= data_in(19);
	wire_w_data_in_range99w(0) <= data_in(1);
	wire_w_data_in_range175w(0) <= data_in(20);
	wire_w_data_in_range179w(0) <= data_in(21);
	wire_w_data_in_range103w(0) <= data_in(2);
	wire_w_data_in_range107w(0) <= data_in(3);
	wire_w_data_in_range111w(0) <= data_in(4);
	wire_w_data_in_range115w(0) <= data_in(5);
	wire_w_data_in_range119w(0) <= data_in(6);
	wire_w_data_in_range123w(0) <= data_in(7);
	wire_w_data_in_range127w(0) <= data_in(8);
	wire_w_data_in_range131w(0) <= data_in(9);
	wire_w_param_decoder_param_latch_range794w(0) <= param_decoder_param_latch(0);
	wire_w_param_decoder_param_latch_range796w(0) <= param_decoder_param_latch(1);
	wire_w_param_decoder_param_latch_range799w(0) <= param_decoder_param_latch(2);
	wire_w_param_decoder_param_latch_range802w(0) <= param_decoder_param_latch(3);
	wire_w_param_decoder_param_latch_range805w(0) <= param_decoder_param_latch(4);
	wire_w_param_decoder_param_latch_range808w(0) <= param_decoder_param_latch(5);
	wire_w_param_decoder_param_latch_range811w(0) <= param_decoder_param_latch(6);
	wire_w_read_source_range1034w(0) <= read_source(0);
	wire_w_read_source_range1038w(0) <= read_source(1);
	wire_w_rsource_parallel_in_range4w(0) <= rsource_parallel_in(0);
	wire_w_rsource_state_par_ini_range12w(0) <= rsource_state_par_ini(0);
	wire_w_rsource_state_par_ini_range16w(0) <= rsource_state_par_ini(1);
	wire_w_wsource_state_par_ini_range22w(0) <= wsource_state_par_ini(0);
	wire_w_wsource_state_par_ini_range26w(0) <= wsource_state_par_ini(1);
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe10 <= (idle AND read_param);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe11 <= ((read_init OR read_source_update) AND wire_w_lg_rsource_update_done957w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe12 <= rsource_update_done;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe13 <= (wire_w_lg_read_init_counter962w(0) OR wire_w_lg_read_pre_data961w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe14 <= (((read_init_counter AND bit_counter_param_start_match) OR (read_pre_data AND bit_counter_param_start_match)) OR (wire_w_lg_read_data966w(0) AND wire_w_lg_width_counter_all_done964w(0)));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe15 <= (((read_data AND width_counter_param_width_match) AND wire_w_lg_width_counter_all_done964w(0)) OR wire_w_lg_read_post972w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe16 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe16 <= (idle AND write_param);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe17 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe17 <= ((write_init OR write_source_update) AND wire_w_lg_wsource_update_done977w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe18 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe18 <= wsource_update_done;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe19 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe19 <= (wire_w_lg_write_init_counter981w(0) OR wire_w_lg_write_pre_data980w(0));
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe1a_ena(0) = '1') THEN dffe1a0 <= (wire_w_lg_rsource_load7w(0) OR wire_w_lg_w_lg_rsource_load5w6w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe1a_ena(1) = '1') THEN dffe1a1 <= (rsource_parallel_in(1) AND rsource_load);
			END IF;
		END IF;
	END PROCESS;
	loop0 : FOR i IN 0 TO 1 GENERATE
		wire_dffe1a_ena(i) <= wire_w_lg_rsource_load1w(0);
	END GENERATE loop0;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe20 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe20 <= (((write_init_counter AND bit_counter_param_start_match) OR (write_pre_data AND bit_counter_param_start_match)) OR (wire_w_lg_write_data984w(0) AND wire_w_lg_bit_counter_all_done983w(0)));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe21 <= (((write_data AND width_counter_param_width_match) AND wire_w_lg_bit_counter_all_done983w(0)) OR wire_w_lg_write_post_data990w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe22 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe22 <= ((write_data AND bit_counter_all_done) OR (write_post_data AND bit_counter_all_done));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe23 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe23 <= write_load;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe24 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe24 <= rublock_regout;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe25a(0) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe25a_ena(0) = '1') THEN dffe25a(0) <= combine_port(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe25a(1) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe25a_ena(1) = '1') THEN dffe25a(1) <= combine_port(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe25a(2) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe25a_ena(2) = '1') THEN dffe25a(2) <= combine_port(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe25a(3) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe25a_ena(3) = '1') THEN dffe25a(3) <= combine_port(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe25a(4) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe25a_ena(4) = '1') THEN dffe25a(4) <= combine_port(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe25a(5) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe25a_ena(5) = '1') THEN dffe25a(5) <= combine_port(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe25a(6) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe25a_ena(6) = '1') THEN dffe25a(6) <= combine_port(6);
			END IF;
		END IF;
	END PROCESS;
	loop1 : FOR i IN 0 TO 6 GENERATE
		wire_dffe25a_ena(i) <= (idle AND (write_param OR read_param));
	END GENERATE loop1;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe2a_ena(0) = '1') THEN dffe2a0 <= (wire_w_lg_rsource_load14w(0) OR wire_w_lg_w_lg_rsource_load5w13w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe2a_ena(1) = '1') THEN dffe2a1 <= (wire_w_lg_rsource_load18w(0) OR wire_w_lg_w_lg_rsource_load5w17w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe2a_ena(2) = '1') THEN dffe2a2 <= (rsource_state_par_ini(2) AND rsource_load);
			END IF;
		END IF;
	END PROCESS;
	loop2 : FOR i IN 0 TO 2 GENERATE
		wire_dffe2a_ena(i) <= wire_w_lg_rsource_load9w(0);
	END GENERATE loop2;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe3a_ena(0) = '1') THEN dffe3a0 <= (wire_w_lg_rsource_load24w(0) OR wire_w_lg_w_lg_rsource_load5w23w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe3a_ena(1) = '1') THEN dffe3a1 <= (wire_w_lg_rsource_load28w(0) OR wire_w_lg_w_lg_rsource_load5w27w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock)
	BEGIN
		IF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe3a_ena(2) = '1') THEN dffe3a2 <= (wsource_state_par_ini(2) AND rsource_load);
			END IF;
		END IF;
	END PROCESS;
	loop3 : FOR i IN 0 TO 2 GENERATE
		wire_dffe3a_ena(i) <= wire_w_lg_rsource_load9w(0);
	END GENERATE loop3;
	PROCESS (clock, wire_dffe7a_clrn(0))
	BEGIN
		IF (wire_dffe7a_clrn(0) = '0') THEN dffe7a(0) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(0) = '1') THEN dffe7a(0) <= (wire_w_lg_shift_reg_load_enable97w(0) OR wire_w_lg_w_lg_shift_reg_load_enable93w96w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(1))
	BEGIN
		IF (wire_dffe7a_clrn(1) = '0') THEN dffe7a(1) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(1) = '1') THEN dffe7a(1) <= (wire_w_lg_shift_reg_load_enable101w(0) OR wire_w_lg_w_lg_shift_reg_load_enable93w100w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(2))
	BEGIN
		IF (wire_dffe7a_clrn(2) = '0') THEN dffe7a(2) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(2) = '1') THEN dffe7a(2) <= (wire_w_lg_shift_reg_load_enable105w(0) OR wire_w_lg_w_lg_shift_reg_load_enable93w104w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(3))
	BEGIN
		IF (wire_dffe7a_clrn(3) = '0') THEN dffe7a(3) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(3) = '1') THEN dffe7a(3) <= (wire_w_lg_shift_reg_load_enable109w(0) OR wire_w_lg_w_lg_shift_reg_load_enable93w108w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(4))
	BEGIN
		IF (wire_dffe7a_clrn(4) = '0') THEN dffe7a(4) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(4) = '1') THEN dffe7a(4) <= (wire_w_lg_shift_reg_load_enable113w(0) OR wire_w_lg_w_lg_shift_reg_load_enable93w112w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(5))
	BEGIN
		IF (wire_dffe7a_clrn(5) = '0') THEN dffe7a(5) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(5) = '1') THEN dffe7a(5) <= (wire_w_lg_shift_reg_load_enable117w(0) OR wire_w_lg_w_lg_shift_reg_load_enable93w116w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(6))
	BEGIN
		IF (wire_dffe7a_clrn(6) = '0') THEN dffe7a(6) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(6) = '1') THEN dffe7a(6) <= (wire_w_lg_shift_reg_load_enable121w(0) OR wire_w_lg_w_lg_shift_reg_load_enable93w120w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(7))
	BEGIN
		IF (wire_dffe7a_clrn(7) = '0') THEN dffe7a(7) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(7) = '1') THEN dffe7a(7) <= (wire_w_lg_shift_reg_load_enable125w(0) OR wire_w_lg_w_lg_shift_reg_load_enable93w124w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(8))
	BEGIN
		IF (wire_dffe7a_clrn(8) = '0') THEN dffe7a(8) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(8) = '1') THEN dffe7a(8) <= (wire_w_lg_shift_reg_load_enable129w(0) OR wire_w_lg_w_lg_shift_reg_load_enable93w128w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(9))
	BEGIN
		IF (wire_dffe7a_clrn(9) = '0') THEN dffe7a(9) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(9) = '1') THEN dffe7a(9) <= (wire_w_lg_shift_reg_load_enable133w(0) OR wire_w_lg_w_lg_shift_reg_load_enable93w132w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(10))
	BEGIN
		IF (wire_dffe7a_clrn(10) = '0') THEN dffe7a(10) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(10) = '1') THEN dffe7a(10) <= (wire_w_lg_shift_reg_load_enable137w(0) OR wire_w_lg_w_lg_shift_reg_load_enable93w136w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(11))
	BEGIN
		IF (wire_dffe7a_clrn(11) = '0') THEN dffe7a(11) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(11) = '1') THEN dffe7a(11) <= (wire_w_lg_shift_reg_load_enable141w(0) OR wire_w_lg_w_lg_shift_reg_load_enable93w140w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(12))
	BEGIN
		IF (wire_dffe7a_clrn(12) = '0') THEN dffe7a(12) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(12) = '1') THEN dffe7a(12) <= (wire_w_lg_shift_reg_load_enable145w(0) OR wire_w_lg_w_lg_shift_reg_load_enable93w144w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(13))
	BEGIN
		IF (wire_dffe7a_clrn(13) = '0') THEN dffe7a(13) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(13) = '1') THEN dffe7a(13) <= (wire_w_lg_shift_reg_load_enable149w(0) OR wire_w_lg_w_lg_shift_reg_load_enable93w148w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(14))
	BEGIN
		IF (wire_dffe7a_clrn(14) = '0') THEN dffe7a(14) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(14) = '1') THEN dffe7a(14) <= (wire_w_lg_shift_reg_load_enable153w(0) OR wire_w_lg_w_lg_shift_reg_load_enable93w152w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(15))
	BEGIN
		IF (wire_dffe7a_clrn(15) = '0') THEN dffe7a(15) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(15) = '1') THEN dffe7a(15) <= (wire_w_lg_shift_reg_load_enable157w(0) OR wire_w_lg_w_lg_shift_reg_load_enable93w156w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(16))
	BEGIN
		IF (wire_dffe7a_clrn(16) = '0') THEN dffe7a(16) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(16) = '1') THEN dffe7a(16) <= (wire_w_lg_shift_reg_load_enable161w(0) OR wire_w_lg_w_lg_shift_reg_load_enable93w160w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(17))
	BEGIN
		IF (wire_dffe7a_clrn(17) = '0') THEN dffe7a(17) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(17) = '1') THEN dffe7a(17) <= (wire_w_lg_shift_reg_load_enable165w(0) OR wire_w_lg_w_lg_shift_reg_load_enable93w164w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(18))
	BEGIN
		IF (wire_dffe7a_clrn(18) = '0') THEN dffe7a(18) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(18) = '1') THEN dffe7a(18) <= (wire_w_lg_shift_reg_load_enable169w(0) OR wire_w_lg_w_lg_shift_reg_load_enable93w168w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(19))
	BEGIN
		IF (wire_dffe7a_clrn(19) = '0') THEN dffe7a(19) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(19) = '1') THEN dffe7a(19) <= (wire_w_lg_shift_reg_load_enable173w(0) OR wire_w_lg_w_lg_shift_reg_load_enable93w172w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(20))
	BEGIN
		IF (wire_dffe7a_clrn(20) = '0') THEN dffe7a(20) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(20) = '1') THEN dffe7a(20) <= (wire_w_lg_shift_reg_load_enable177w(0) OR wire_w_lg_w_lg_shift_reg_load_enable93w176w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(21))
	BEGIN
		IF (wire_dffe7a_clrn(21) = '0') THEN dffe7a(21) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(21) = '1') THEN dffe7a(21) <= (wire_w_lg_shift_reg_load_enable181w(0) OR wire_w_lg_w_lg_shift_reg_load_enable93w180w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(22))
	BEGIN
		IF (wire_dffe7a_clrn(22) = '0') THEN dffe7a(22) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(22) = '1') THEN dffe7a(22) <= (wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(23));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(23))
	BEGIN
		IF (wire_dffe7a_clrn(23) = '0') THEN dffe7a(23) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(23) = '1') THEN dffe7a(23) <= (wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(24));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(24))
	BEGIN
		IF (wire_dffe7a_clrn(24) = '0') THEN dffe7a(24) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(24) = '1') THEN dffe7a(24) <= (wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(25));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(25))
	BEGIN
		IF (wire_dffe7a_clrn(25) = '0') THEN dffe7a(25) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(25) = '1') THEN dffe7a(25) <= (wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(26));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(26))
	BEGIN
		IF (wire_dffe7a_clrn(26) = '0') THEN dffe7a(26) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(26) = '1') THEN dffe7a(26) <= (wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(27));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(27))
	BEGIN
		IF (wire_dffe7a_clrn(27) = '0') THEN dffe7a(27) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(27) = '1') THEN dffe7a(27) <= (wire_w_lg_shift_reg_load_enable93w(0) AND dffe7a(28));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe7a_clrn(28))
	BEGIN
		IF (wire_dffe7a_clrn(28) = '0') THEN dffe7a(28) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe7a_ena(28) = '1') THEN dffe7a(28) <= (wire_w_lg_shift_reg_load_enable93w(0) AND shift_reg_serial_in);
			END IF;
		END IF;
	END PROCESS;
	loop4 : FOR i IN 0 TO 28 GENERATE
		wire_dffe7a_clrn(i) <= wire_w_lg_w_lg_shift_reg_clear91w92w(0);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 28 GENERATE
		wire_dffe7a_ena(i) <= wire_w_lg_shift_reg_load_enable90w(0);
	END GENERATE loop5;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe8 <= '1';
		ELSIF (clock = '1' AND clock'event) THEN dffe8 <= (((wire_w_lg_w_lg_w_lg_idle949w950w951w(0) OR (read_data AND width_counter_all_done)) OR (read_post AND width_counter_all_done)) OR power_up);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe9 <= ((((wire_w_lg_w_lg_w_lg_idle949w950w951w(0) OR (read_data AND width_counter_all_done)) OR (read_post AND width_counter_all_done)) OR power_up) AND write_load);
		END IF;
	END PROCESS;
	wire_cntr5_w_lg_w_q_range30w33w(0) <= wire_cntr5_w_q_range30w(0) AND wire_cntr5_w_lg_w_q_range31w32w(0);
	wire_cntr5_w_lg_w_q_range31w32w(0) <= NOT wire_cntr5_w_q_range31w(0);
	wire_cntr5_w_q_range30w(0) <= wire_cntr5_q(0);
	wire_cntr5_w_q_range31w(0) <= wire_cntr5_q(1);
	cntr5 :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 6
	  )
	  PORT MAP ( 
		clock => clock,
		cnt_en => bit_counter_enable,
		q => wire_cntr5_q,
		sclr => bit_counter_clear
	  );
	cntr6 :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 5
	  )
	  PORT MAP ( 
		clock => clock,
		cnt_en => width_counter_enable,
		q => wire_cntr6_q,
		sclr => width_counter_clear
	  );
	sd4 :  cycloneive_rublock
	  PORT MAP ( 
		captnupdt => rublock_captnupdt,
		clk => rublock_clock,
		rconfig => rublock_reconfig,
		regin => rublock_regin,
		regout => wire_sd4_regout,
		rsttimer => reset_timer,
		shiftnld => rublock_shiftnld
	  );

 END RTL; --altremote_rmtupdt_51n
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY altremote IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		data_in		: IN STD_LOGIC_VECTOR (21 DOWNTO 0);
		param		: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		read_param		: IN STD_LOGIC ;
		read_source		: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
		reconfig		: IN STD_LOGIC ;
		reset		: IN STD_LOGIC ;
		reset_timer		: IN STD_LOGIC ;
		write_param		: IN STD_LOGIC ;
		busy		: OUT STD_LOGIC ;
		data_out		: OUT STD_LOGIC_VECTOR (28 DOWNTO 0)
	);
END altremote;


ARCHITECTURE RTL OF altremote IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "altremote_update";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "check_app_pof=false;intended_device_family=Cyclone IV E;in_data_width=22;operation_mode=REMOTE;out_data_width=29;";
	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (28 DOWNTO 0);



	COMPONENT altremote_rmtupdt_51n
	PORT (
			clock	: IN STD_LOGIC ;
			data_in	: IN STD_LOGIC_VECTOR (21 DOWNTO 0);
			read_param	: IN STD_LOGIC ;
			read_source	: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
			busy	: OUT STD_LOGIC ;
			data_out	: OUT STD_LOGIC_VECTOR (28 DOWNTO 0);
			param	: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			reconfig	: IN STD_LOGIC ;
			reset	: IN STD_LOGIC ;
			reset_timer	: IN STD_LOGIC ;
			write_param	: IN STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	busy    <= sub_wire0;
	data_out    <= sub_wire1(28 DOWNTO 0);

	altremote_rmtupdt_51n_component : altremote_rmtupdt_51n
	PORT MAP (
		clock => clock,
		data_in => data_in,
		read_param => read_param,
		read_source => read_source,
		param => param,
		reconfig => reconfig,
		reset => reset,
		reset_timer => reset_timer,
		write_param => write_param,
		busy => sub_wire0,
		data_out => sub_wire1
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: PRIVATE: SIM_INIT_CONFIG_COMBO STRING "FACTORY"
-- Retrieval info: PRIVATE: SIM_INIT_PAGE_SELECT_COMBO STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT0_CHECK STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT1_CHECK STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT2_CHECK STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT3_CHECK STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT4_CHECK STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_WATCHDOG_VALUE_EDIT STRING "1"
-- Retrieval info: PRIVATE: SUPPORT_WRITE_CHECK STRING "1"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: WATCHDOG_ENABLE_CHECK STRING "0"
-- Retrieval info: CONSTANT: CHECK_APP_POF STRING "false"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: IN_DATA_WIDTH NUMERIC "22"
-- Retrieval info: CONSTANT: OPERATION_MODE STRING "REMOTE"
-- Retrieval info: CONSTANT: OUT_DATA_WIDTH NUMERIC "29"
-- Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: data_in 0 0 22 0 INPUT NODEFVAL "data_in[21..0]"
-- Retrieval info: USED_PORT: data_out 0 0 29 0 OUTPUT NODEFVAL "data_out[28..0]"
-- Retrieval info: USED_PORT: param 0 0 3 0 INPUT NODEFVAL "param[2..0]"
-- Retrieval info: USED_PORT: read_param 0 0 0 0 INPUT NODEFVAL "read_param"
-- Retrieval info: USED_PORT: read_source 0 0 2 0 INPUT NODEFVAL "read_source[1..0]"
-- Retrieval info: USED_PORT: reconfig 0 0 0 0 INPUT NODEFVAL "reconfig"
-- Retrieval info: USED_PORT: reset 0 0 0 0 INPUT NODEFVAL "reset"
-- Retrieval info: USED_PORT: reset_timer 0 0 0 0 INPUT NODEFVAL "reset_timer"
-- Retrieval info: USED_PORT: write_param 0 0 0 0 INPUT NODEFVAL "write_param"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @data_in 0 0 22 0 data_in 0 0 22 0
-- Retrieval info: CONNECT: @param 0 0 3 0 param 0 0 3 0
-- Retrieval info: CONNECT: @read_param 0 0 0 0 read_param 0 0 0 0
-- Retrieval info: CONNECT: @read_source 0 0 2 0 read_source 0 0 2 0
-- Retrieval info: CONNECT: @reconfig 0 0 0 0 reconfig 0 0 0 0
-- Retrieval info: CONNECT: @reset 0 0 0 0 reset 0 0 0 0
-- Retrieval info: CONNECT: @reset_timer 0 0 0 0 reset_timer 0 0 0 0
-- Retrieval info: CONNECT: @write_param 0 0 0 0 write_param 0 0 0 0
-- Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
-- Retrieval info: CONNECT: data_out 0 0 29 0 @data_out 0 0 29 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL altremote.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altremote.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altremote.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altremote.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altremote_inst.vhd TRUE
-- Retrieval info: LIB_FILE: cycloneive
-- Retrieval info: LIB_FILE: lpm
