altremote_inst : altremote PORT MAP (
		clock	 => clock_sig,
		data_in	 => data_in_sig,
		param	 => param_sig,
		read_param	 => read_param_sig,
		read_source	 => read_source_sig,
		reconfig	 => reconfig_sig,
		reset	 => reset_sig,
		reset_timer	 => reset_timer_sig,
		write_param	 => write_param_sig,
		busy	 => busy_sig,
		data_out	 => data_out_sig
	);
